module pc_module #(
    parameter DATA_WIDTH = 32
) (
    input  logic                    clk,
    input  logic                    rst,
    input  logic [DATA_WIDTH-1:0]   PCNext_i,
    output logic [DATA_WIDTH-1:0]   PC_o
);

    logic [DATA_WIDTH-1:0] PC;

    always_ff @(posedge clk) begin
        if (rst) 
            PC <= {DATA_WIDTH{1'b0}};
        else 
            PC <= PCNext_i;
    end

    always_comb begin
        PC_o = PC;
    end

endmodule
